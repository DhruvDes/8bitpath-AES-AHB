`include "ahb_if.svh"

package ahb_pkg;

`include "uvm_macros.svh"
import uvm_pkg :: *;



`include "ahb_common.sv"
`include "ahb_tx.sv"
`include "ahb_seq_lib.sv"
// // `include "ahb_sqr.sv"
`include "ahb_drv.sv"
`include "ahb_mon.sv"
`include "ahb_cov.sv"
`include "ahb_agent_m.sv"
`include "ahb_env.sv"
`include "test_lib.sv" 


endpackage