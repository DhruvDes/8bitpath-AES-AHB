package master_agent_pkg;


`include "uvm_macros.svh"
import uvm_pkg :: *;

`include "common.sv"
`include "m_a_trnsaction.sv"











endpackage