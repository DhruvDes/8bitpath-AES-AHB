package aes_pkg;

 
  import uvm_pkg::*;
  `include "uvm_macros.svh"



  `include "tran.sv"          
  `include "monitor.sv"       
  `include "driver.sv"        
  `include "agnt.sv"          
  `include "scrbrd.sv"        
  `include "envr.sv"          
  `include "seq_library.sv"   
  `include "test.sv"          

endpackage : aes_pkg
