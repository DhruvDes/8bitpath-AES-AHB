package ahb_pkg;

`include "uvm_macros.svh"
import uvm_pkg :: *;

`include "ahb_interface.sv"
import interfaces :: *;

`include "ahb_common.sv"
`include "ahb_tx.sv"
`include "ahb_seq_lib.sv"
// `include "ahb_sqr.sv"
`include "ahb_drv.sv"
`include "ahb_agent.sv"
`include "ahb_env.sv"
`include "test_lib.sv" 


endpackage