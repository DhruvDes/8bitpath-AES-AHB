
package ahb_pkg;
`include "uvm_macros.svh"
import uvm_pkg :: *;


`include "ahb_trn.sv"
`include "ahb_seq_lib.sv"

// // `include "ahb_sqr.sv"
`include "ahb_drv.sv"
`include "ahb_mon.sv"
`include "ahb_scb.sv"
`include "ahb_cover.sv"
`include "ahb_agent.sv"
`include "ahb_subor.sv"
`include "sub_agent.sv"
`include "ahb_env.sv"
`include "test_lib.sv" 


endpackage